library verilog;
use verilog.vl_types.all;
entity Crossbar_vlg_tst is
    generic(
        count           : integer := 2
    );
end Crossbar_vlg_tst;
