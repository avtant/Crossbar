library verilog;
use verilog.vl_types.all;
entity Crossbar_vlg_tst is
end Crossbar_vlg_tst;
